//non